-- A DUT entity is used to wrap your design so that we can combine it with testbench.
-- This example shows how you can do this for the OR Gate

library ieee;
use ieee.std_logic_1164.all;

entity DUT is
    port(input_vector: in std_logic_vector(2 downto 0);
       	output_vector: out std_logic_vector(2 downto 0));
end entity;

architecture DutWrap of DUT is
   component seq_gen is
     port(UD, reset, clock: in std_logic; y: out std_logic_vector);
   end component;
begin

   -- input/output vector element ordering is critical,
   -- and must match the ordering in the trace file!
   add_instance: seq_gen
			port map (
					UD => input_vector(2),
					reset => input_vector(1),
					clock => input_vector(0),
					y => output_vector(2 downto 0));
end DutWrap;